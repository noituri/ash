main =
//    log.info "test" <- Logger that needs to be implemented
    println "test"