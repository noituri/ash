main =
//    log.info "test" <- Logger that needs to be implemented */
    println /* comment test */ "123"
    println(321)