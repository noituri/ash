main =>
    test
    test2
    ff(a, b)(aaaaa,bbb)
    ff -12, b(-14.23), 32
    ff (a), b, c, aa bb, cc
    // comment test
    // println /* comment test 2 */ "test"
    // println(123)
