main =>
    test
    test2
        ff
                
    // comment test
    // println /* comment test 2 */ "test"
    // println(123)