main =>
    test
    test2
    ff(a, b)(aaaaa,bbb)
    ff a, b                
    // comment test
    // println /* comment test 2 */ "test"
    // println(123)