main =>
    test
    test2
    ff(a, b)(aaaaa,bbb)
    // comment test
    // println /* comment test 2 */ "test"
    // println(123)